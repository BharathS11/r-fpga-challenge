// /r/fpga challenge
//
// This is the interface for the component for this week
// It's a counter; it should reset to 0 when `reset` is driven to 1
// and count up when `enable` is driven to 1
module challenge(input clk, input reset, input enable, output [3:0] count);
// TODO: some code!
endmodule
